	0 => X"61",
	1 => X"00",
	2 => X"00",
	3 => X"61",
	4 => X"01",
	5 => X"03",
	6 => X"61",
	7 => X"02",
	8 => X"02",
	9 => X"69",
	10 => X"02",
	11 => X"00",
	12 => X"6d",
	13 => X"16",
	14 => X"63",
	15 => X"02",
	16 => X"01",
	17 => X"02",
	18 => X"00",
	19 => X"01",
	20 => X"67",
	21 => X"09",
	22 => X"61",
	23 => X"03",
	24 => X"01",
	25 => X"61",
	26 => X"01",
	27 => X"02",
	28 => X"01",
	29 => X"02",
	30 => X"00",
	31 => X"69",
	32 => X"02",
	33 => X"00",
	34 => X"6d",
	35 => X"3f",
	36 => X"61",
	37 => X"04",
	38 => X"00",
	39 => X"61",
	40 => X"05",
	41 => X"02",
	42 => X"69",
	43 => X"05",
	44 => X"00",
	45 => X"6d",
	46 => X"37",
	47 => X"02",
	48 => X"04",
	49 => X"03",
	50 => X"63",
	51 => X"05",
	52 => X"01",
	53 => X"67",
	54 => X"2a",
	55 => X"01",
	56 => X"03",
	57 => X"04",
	58 => X"63",
	59 => X"02",
	60 => X"01",
	61 => X"67",
	62 => X"1f",
	63 => X"08",
	64 => X"03",
	65 => X"00",
