	0 => X"28",
	1 => X"03",
